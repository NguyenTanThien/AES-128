library verilog;
use verilog.vl_types.all;
entity InvMixColumns is
    port(
        \IN\            : in     vl_logic_vector(127 downto 0);
        \OUT\           : out    vl_logic_vector(127 downto 0)
    );
end InvMixColumns;
