library verilog;
use verilog.vl_types.all;
entity ShiftRows is
    port(
        s               : in     vl_logic_vector(127 downto 0);
        s1              : out    vl_logic_vector(127 downto 0)
    );
end ShiftRows;
